module dont_kill_top_level (
	input clk,    // Clock
	input resetn, //active low reset
	
);

  

endmodule

